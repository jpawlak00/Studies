`timescale 1ns / 1ps
module char_rom_16x16(
  output reg [6:0] char_code,
  
  input wire [7:0] char_xy
  );
  
 always @*
         case (char_xy)
             //code x00
             8'h00: char_code = 7'h0c;
             8'h01: char_code = 7'h0c;
             8'h02: char_code = 7'h0c;
             8'h03: char_code = 7'h0c;
             8'h04: char_code = 7'h0c;
             8'h05: char_code = 7'h0c;
             8'h06: char_code = 7'h0c;
             8'h07: char_code = 7'h0c;
             8'h08: char_code = 7'h0c;
             8'h09: char_code = 7'h0c;
             8'h0a: char_code = 7'h0c;
             8'h0b: char_code = 7'h0c;
             8'h0c: char_code = 7'h0c;
             8'h0d: char_code = 7'h0c;
             8'h0e: char_code = 7'h0c;
             8'h0f: char_code = 7'h0c;
             8'h10: char_code = 7'h0c;
             8'h11: char_code = 7'h0c;
             8'h12: char_code = 7'h0c;
             8'h13: char_code = 7'h0c;
             8'h14: char_code = 7'h0c;
             8'h15: char_code = 7'h0c;
             8'h16: char_code = 7'h0c;
             8'h17: char_code = 7'h0c;
             8'h18: char_code = 7'h0c;
             8'h19: char_code = 7'h0c;
             8'h1a: char_code = 7'h0c;
             8'h1b: char_code = 7'h0c;
             8'h1c: char_code = 7'h0c;
             8'h1d: char_code = 7'h0c;
             8'h1e: char_code = 7'h0c;
             8'h1f: char_code = 7'h0c;
             8'h20: char_code = 7'h0c;
             8'h21: char_code = 7'h0c;
             8'h22: char_code = 7'h0c;
             8'h23: char_code = 7'h0c;
             8'h24: char_code = 7'h0c;
             8'h25: char_code = 7'h0c;
             8'h26: char_code = 7'h0c;
             8'h27: char_code = 7'h0c;
             8'h28: char_code = 7'h0c;
             8'h29: char_code = 7'h0c;
             8'h2a: char_code = 7'h0c;
             8'h2b: char_code = 7'h0c;
             8'h2c: char_code = 7'h0c;
             8'h2d: char_code = 7'h0c;
             8'h2e: char_code = 7'h0c;
             8'h2f: char_code = 7'h0c;
             8'h30: char_code = 7'h0c;
             8'h31: char_code = 7'h0c;
             8'h32: char_code = 7'h0c;
             8'h33: char_code = 7'h0c;
             8'h34: char_code = 7'h0c;
             8'h35: char_code = 7'h0c;
             8'h36: char_code = 7'h0c;
             8'h37: char_code = 7'h0c;
             8'h38: char_code = 7'h0c;
             8'h39: char_code = 7'h0c;
             8'h3a: char_code = 7'h0c;
             8'h3b: char_code = 7'h0c;
             8'h3c: char_code = 7'h0c;
             8'h3d: char_code = 7'h0c;
             8'h3e: char_code = 7'h0c;
             8'h3f: char_code = 7'h0c;
             8'h40: char_code = 7'h0c;
             8'h41: char_code = 7'h0c;
             8'h42: char_code = 7'h0c;
             8'h43: char_code = 7'h0c;
             8'h44: char_code = 7'h0c;
             8'h45: char_code = 7'h0c;
             8'h46: char_code = 7'h0c;
             8'h47: char_code = 7'h0c;
             8'h48: char_code = 7'h0c;
             8'h49: char_code = 7'h0c;
             8'h4a: char_code = 7'h0c;
             8'h4b: char_code = 7'h0c;
             8'h4c: char_code = 7'h0c;
             8'h4d: char_code = 7'h0c;
             8'h4e: char_code = 7'h0c;
             8'h4f: char_code = 7'h0c;
             8'h50: char_code = 7'h0c;
             8'h51: char_code = 7'h0c;
             8'h52: char_code = 7'h0c;
             8'h53: char_code = 7'h0c;
             8'h54: char_code = 7'h0c;
             8'h55: char_code = 7'h0c;
             8'h56: char_code = 7'h0c;
             8'h57: char_code = 7'h0c;
             8'h58: char_code = 7'h0c;
             8'h59: char_code = 7'h0c;
             8'h5a: char_code = 7'h0c;
             8'h5b: char_code = 7'h0c;
             8'h5c: char_code = 7'h0c;
             8'h5d: char_code = 7'h0c;
             8'h5e: char_code = 7'h0c;
             8'h5f: char_code = 7'h0c;
             8'h60: char_code = 7'h0c;
             8'h61: char_code = 7'h0c;
             8'h62: char_code = 7'h0c;
             8'h63: char_code = 7'h0c;
             8'h64: char_code = 7'h0c;
             8'h65: char_code = 7'h0c;
             8'h66: char_code = 7'h0c;
             8'h67: char_code = 7'h0c;
             8'h68: char_code = 7'h0c;
             8'h69: char_code = 7'h0c;
             8'h6a: char_code = 7'h0c;
             8'h6b: char_code = 7'h0c;
             8'h6c: char_code = 7'h0c;
             8'h6d: char_code = 7'h0c;
             8'h6e: char_code = 7'h0c;
             8'h6f: char_code = 7'h0c;
             8'h70: char_code = 7'h0c;
             8'h71: char_code = 7'h0c;
             8'h72: char_code = 7'h0c;
             8'h73: char_code = 7'h0c;
             8'h74: char_code = 7'h0c;
             8'h75: char_code = 7'h0c;
             8'h76: char_code = 7'h0c;
             8'h77: char_code = 7'h0c;
             8'h78: char_code = 7'h0c;
             8'h79: char_code = 7'h0c;
             8'h7a: char_code = 7'h0c;
             8'h7b: char_code = 7'h0c;
             8'h7c: char_code = 7'h0c;
             8'h7d: char_code = 7'h0c;
             8'h7e: char_code = 7'h0c;
             8'h7f: char_code = 7'h0c;
        endcase
endmodule
